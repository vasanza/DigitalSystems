library ieee;
use ieee.std_logic_1164.all;

entity ContUp is
	port(resetn,en,clk: in std_logic;
				Qout: out std_logic_vector(3 downto 0));
end ContUp;

architecture comp of ContUp is
		begin
end comp;