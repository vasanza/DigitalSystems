LIBRARY IEEE;
USE  IEEE.STD_LOGIC_1164.all;
USE  IEEE.STD_LOGIC_UNSIGNED.all;

ENTITY Comp IS
	Port(A,B : in std_logic_vector(3 downto 0);
			AmayB,AmenB : out std_logic);
END Comp;

ARCHITECTURE sol OF Comp IS
BEGIN

END sol;