library ieee;
use ieee.std_logic_1164.all;

entity RAM is
	port(Add,Din: in std_logic_vector(3 downto 0);
				clk,modo: in std_logic;
				Dout: out std_logic_vector(3 downto 0));
end RAM;

architecture comp of RAM is
		begin
end comp;