library ieee;
use ieee.std_logic_1164.all;

entity MSS is
	port(restn,st,fin,clk: in std_logic;
				ResetCnt,ecnt,ei,et,edeco: out std_logic);
end MSS;

architecture comp of MSS is
		begin
end comp;