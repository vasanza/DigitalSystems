library ieee;
use ieee.std_logic_1164.all;

entity RegAcum is
	port(Din: in std_logic_vector(3 downto 0);
				clk,en: in std_logic;
				Qout: out std_logic_vector(3 downto 0));
end RegAcum;

architecture comp of RegAcum is
		begin
end comp;