library ieee;
use ieee.std_logic_1164.all;

Entity mss is
	Port(	AmaB,AmeB,Resetn,Clk,Start,KeyIn,FinCnt: in std_logic;
			eDeco,m,eMin,eMax,modo,eCnt,ResetnCnt: out std_logic);
end mss;

Architecture sol of mss is
Begin

end sol;