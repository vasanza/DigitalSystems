LIBRARY IEEE;
USE  IEEE.STD_LOGIC_1164.all;
USE  IEEE.STD_LOGIC_UNSIGNED.all;

ENTITY KeyDeco IS
	Port(Key : in std_logic_vector(3 downto 0);
			Q : out std_logic_vector(3 downto 0));
END KeyDeco;

ARCHITECTURE sol OF KeyDeco IS
BEGIN

END sol;