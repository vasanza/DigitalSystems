library ieee;
use ieee.std_logic_1164.all;

entity MUX is
	port(D0,D1: in std_logic_vector(3 downto 0);
				m: in std_logic;
				Qout: out std_logic_vector(3 downto 0));
end MUX;

architecture comp of MUX is
		begin
end comp;