library ieee;
use ieee.std_logic_1164.all;

entity DecoInst is
	port(Din: in std_logic_vector(3 downto 0);
				en,clk: in std_logic;
				fin,modo,m,s,ea: out std_logic);
end DecoInst;

architecture comp of DecoInst is
		begin
end comp;