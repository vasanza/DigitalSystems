library ieee;
use ieee.std_logic_1164.all;

entity ALU is
	port(A,B: in std_logic_vector(3 downto 0);
				S: in std_logic;
				Qout: out std_logic_vector(3 downto 0));
end ALU;

architecture comp of ALU is
		begin
end comp;