LIBRARY IEEE;
USE  IEEE.STD_LOGIC_1164.all;
USE  IEEE.STD_LOGIC_UNSIGNED.all;

ENTITY CntUp IS
	Port(en,ResetnCnt,Clk: in std_logic;
			Q : out std_logic_vector(3 downto 0));
END CntUp;

ARCHITECTURE sol OF CntUp IS
BEGIN

END sol;